** Profile: "SCHEMATIC1-Vout"  [ C:\Users\John\Desktop\Elec1\Simulation\Bonus\Part3\vout_full_wave-schematic1-vout.sim ] 

** Creating circuit file "vout_full_wave-schematic1-vout.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80ms 40ms 1us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\vout_full_wave-SCHEMATIC1.net" 


.END
