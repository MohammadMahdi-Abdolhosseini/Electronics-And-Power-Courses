** Profile: "SCHEMATIC1-Part2_Gain"  [ C:\Users\John\Desktop\Elec1\Simulation\Part2\part2-schematic1-part2_gain.sim ] 

** Creating circuit file "part2-schematic1-part2_gain.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0.5ms 1us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part2-SCHEMATIC1.net" 


.END
