** Profile: "SCHEMATIC1-Vout_HALF"  [ C:\USERS\JOHN\DESKTOP\ELEC1\Simulation\Bonus\Part3\bonus_part3-SCHEMATIC1-Vout_HALF.sim ] 

** Creating circuit file "bonus_part3-SCHEMATIC1-Vout_HALF.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.2s 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\bonus_part3-SCHEMATIC1.net" 


.END
