** Profile: "SCHEMATIC1-Vout_FULL"  [ C:\Users\John\Desktop\Elec1\Simulation\Bonus\Part3\vout_full_wave-schematic1-vout_full.sim ] 

** Creating circuit file "vout_full_wave-schematic1-vout_full.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.2s 0 10us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\vout_full_wave-SCHEMATIC1.net" 


.END
