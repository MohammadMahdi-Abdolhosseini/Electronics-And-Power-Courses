** Profile: "SCHEMATIC1-Part1_MaxSwingVCE"  [ C:\Users\John\Desktop\Elec1\Simulation\Part1_CommonCollector\part1_commoncollector-schematic1-part1_maxswingvce.sim ] 

** Creating circuit file "part1_commoncollector-schematic1-part1_maxswingvce.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 10ns 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part1_commoncollector-SCHEMATIC1.net" 


.END
