** Profile: "SCHEMATIC1-Vout_Full_Wave"  [ C:\USERS\JOHN\DESKTOP\ELEC1\Simulation\Bonus\Part2\full_wave_rectifier-SCHEMATIC1-Vout_Full_Wave.sim ] 

** Creating circuit file "full_wave_rectifier-SCHEMATIC1-Vout_Full_Wave.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.1s 0 10us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\full_wave_rectifier-SCHEMATIC1.net" 


.END
