** Profile: "SCHEMATIC1-Vout_HALF_FULL"  [ C:\USERS\JOHN\DESKTOP\ELEC1\Simulation\Bonus\Part2.5\both_wave_rectifier-SCHEMATIC1-Vout_HALF_FULL.sim ] 

** Creating circuit file "both_wave_rectifier-SCHEMATIC1-Vout_HALF_FULL.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.08s 0s 10us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\both_wave_rectifier-SCHEMATIC1.net" 


.END
