** Profile: "SCHEMATIC1-Gain"  [ C:\Users\John\Desktop\Elec1\Simulation\Bonus\Part3\vout_full_wave-SCHEMATIC1-Gain.sim ] 

** Creating circuit file "vout_full_wave-SCHEMATIC1-Gain.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 47ms 46.5ms 1us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\vout_full_wave-SCHEMATIC1.net" 


.END
