** Profile: "SCHEMATIC1-Part2_MaxSwingVEC"  [ C:\Users\John\Desktop\Elec1\Simulation\Part2\part2-SCHEMATIC1-Part2_MaxSwingVEC.sim ] 

** Creating circuit file "part2-SCHEMATIC1-Part2_MaxSwingVEC.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1ms 0 1us 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\part2-SCHEMATIC1.net" 


.END
